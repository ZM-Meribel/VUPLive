<?xml version="1.0" standalone="no"?><!DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd"><svg t="1651276029088" class="icon" viewBox="0 0 1024 1024" version="1.1" xmlns="http://www.w3.org/2000/svg" p-id="6748" xmlns:xlink="http://www.w3.org/1999/xlink" width="200" height="200"><defs><style type="text/css">@font-face { font-family: feedback-iconfont; src: url("//at.alicdn.com/t/font_1031158_u69w8yhxdu.woff2?t=1630033759944") format("woff2"), url("//at.alicdn.com/t/font_1031158_u69w8yhxdu.woff?t=1630033759944") format("woff"), url("//at.alicdn.com/t/font_1031158_u69w8yhxdu.ttf?t=1630033759944") format("truetype"); }
</style></defs><path d="M252.779462 486.963907c11.152909-27.35251 19.517591-55.318431 33.709668-79.994243 22.026996-38.589067 48.124804-74.836022 72.10356-112.33768 8.197388-12.853728 15.530426-26.348748 22.528877-39.927415 5.576455-10.678911 4.070812-18.904181-8.727152-24.369107a155.778262 155.778262 0 0 1-33.793316-19.266651c-9.173268-7.026333-17.482186-7.054215-27.101569-3.234344S292.093467 215.641503 280.940558 216.784677l41.82341-16.729364c-11.152909-15.279486-24.64793-2.481522-37.501658-5.325515L308.822831 188.121699C303.497317 161.968127 278.15233 167.321523 260.502851 155.471557c8.364682-5.855277 15.028545-11.152909 22.305819-15.363133C303.246377 127.812342 314.594462 109.772511 318.916214 86.46293c0.836468-4.516928 4.684222-8.559858 7.444567-12.602787 6.970568-10.316441 15.279486-19.935826 20.883823-30.949324 7.054215-13.941137 6.608099-28.495684-3.9314-42.910819 28.746624 5.855277 48.821861 46.256692 47.037395 92.011503 4.098694-0.557645 7.918566-1.338349 11.738437-1.505643 19.824296-1.003762 39.704358-1.645054 59.528654-2.788227a24.03452 24.03452 0 0 0 12.073025-4.04293c23.588403-17.036069 39.286123-39.035183 43.914581-69.148038 1.728701 6.050453 2.593051 12.519141 5.381278 18.067713 4.461164 8.922328 8.810798 18.625359 15.725603 25.484398 9.20115 9.089621 12.909493 18.597476 11.543261 31.088735-1.003762 9.20115-3.624696 19.517591-0.585528 27.547686s11.40385 15.251604 18.820535 20.995352c7.862801 6.106218 10.037618 11.626908 3.819871 19.684885a180.175252 180.175252 0 0 0-10.874087 14.387253c-1.784466 2.788227-1.979641 6.635981-3.206461 9.898207s-1.895995 7.751272-4.349635 9.31268c-10.595264 6.74751-18.904181 16.06019-29.834032 22.835582-27.240981 16.729364-57.075014 22.8077-87.494575 28.32839a18.430183 18.430183 0 0 0-10.846204 5.269749c-22.556759 29.889797-44.611638 60.560298-41.656117 100.376185 0.97588 12.602788 5.046692 28.216861 13.522903 36.442131 43.998228 42.576232 67.279926 94.79973 77.763661 153.826504 3.541049 20.047355 6.608099 40.150474 10.288559 62.707233 23.337463-1.421996 47.70657-2.788227 72.019912-4.65634 1.979641-0.167294 5.046692-4.29387 5.241868-6.775392 1.561407-18.987828 10.846204-34.546137 21.971231-48.933391 33.737551-43.552111 26.432395-79.380833-11.599026-111.947328a53.980082 53.980082 0 0 1-5.576454-6.74751c10.204912-7.946448 16.729364-1.700819 23.030758 4.377517 35.68931 35.131665 38.477537 79.35295 8.197388 119.44766-7.779154 10.316441-15.753485 20.939587-20.911705 32.650142-5.799513 13.132551-1.505643 17.342774 12.658552 16.729364 9.591502-0.418234 19.238769 0 29.91768 0-6.022571-29.387916 4.489046-51.805264 20.270412-73.051556a109.577335 109.577335 0 0 0 13.745961-25.707457c5.994689-15.502544 4.321752-30.41956-8.22527-42.381055-8.364682-8.002213-18.095596-14.610311-26.209337-22.835582-3.485284-3.513166-4.433281-9.535738-4.321753-15.558309 20.521353 11.822084 40.038945 23.588403 49.992917 45.113519 7.72339 16.729364 5.966807 33.626022-3.206462 49.463153-7.444567 12.825846-15.920778 25.094046-23.225934 38.003539a61.480413 61.480413 0 0 0-7.388802 19.350297c-3.457402 20.605 2.45364 26.376631 23.002875 27.519804 31.953085 1.728701 63.850406 4.823633 95.803492 7.054216 10.288559 0.724939 15.056428 4.238106 12.770082 15.669837-2.788227 13.634432-3.485284 27.631333-5.855278 41.349412-1.394114 8.141624 0 12.491259 8.866563 15.251604 57.716306 17.761008 108.071692 48.738214 154.216855 87.215751 12.519141 10.42797 17.398539 23.198052 17.28701 39.035183-0.223058 38.75636-14.638194 71.350738-41.544588 98.759013C856.737388 939.6605 815.164919 978.528389 763.499066 1003.789729a145.963702 145.963702 0 0 1-93.795968 11.794202c-40.206238-8.085859-80.050007-5.966807-120.451422-0.446116-35.745075 4.879398-72.019913 5.938924-108.099574 7.918565-20.855941 1.115291-41.82341 1.059526-62.679351 0.752822a45.420224 45.420224 0 0 1-18.681124-4.572693A533.527304 533.527304 0 0 1 216.811329 918.497854c-4.600575-4.572693-8.504093-9.842443-12.658552-14.833369C193.334454 890.587699 181.372959 878.319498 172.199691 864.099539c-6.273512-9.535738-13.021022-22.026996-11.989378-32.427084a241.098019 241.098019 0 0 1 15.335251-65.941577c4.405399-10.874087 17.482186-20.103119 28.774506-25.763221 9.870325-4.935162 12.184554-8.225271 10.5395-19.183004-7.305156-48.31998 0.446116-95.998668 14.693958-141.64195 10.567382-33.876962 6.217747-64.129229-7.500332-94.269966A1034.962111 1034.962111 0 0 0 116.435144 301.658317C73.607972 242.938249 79.435367 180.314663 110.579867 118.611192c11.599026-23.030758 53.338789-27.631333 72.493911-9.619385a24.564283 24.564283 0 0 1 6.942686 11.794202c5.911042 27.408275 6.49657 54.649256-7.026333 80.217301-10.344323 19.517591-26.348748 31.534851-49.407389 29.610974-5.576455-0.473999-10.595264-5.994689-15.865013-9.20115 4.684222-3.513166 9.229033-9.703031 14.10843-10.009736 14.164195-0.86435 26.7391-2.537287 33.84908-17.008187 8.364682-17.063951 14.498782-34.155785 7.277273-53.394554s-22.026996-24.926753-38.087185-12.100906a64.352287 64.352287 0 0 0-20.35406 26.962158c-21.525115 60.95065-4.433281 114.066381 32.733789 164.505414 31.674263 42.910819 60.169946 88.191631 89.418451 132.886915 6.74751 10.17703 10.818322 22.250054 16.115955 33.709669z m46.061515 254.119041q3.290108-8.699269 6.635982-17.398539l-2.537287-1.449878-8.531976 7.026333c-8.727152-10.623146-12.296083 3.541049-22.138525 3.568931 21.329939 2.788227 1.533525 9.647267 6.886921 16.729364a66.610751 66.610751 0 0 1 10.901969-8.95021c2.258464-1.198938 5.88316 0.195176 8.894446 0.418235a21.302057 21.302057 0 0 1-2.983404 4.489046c-8.866563 8.225271-9.898207 17.761008-3.178579 27.213099s16.255365 15.112192 27.519804 10.623146 14.275724-15.140075 12.825846-26.543925c-2.397876-18.848417-13.49502-23.727815-34.295197-15.725602z m74.80814-117.997782a26.069926 26.069926 0 0 0-0.975879 5.827396c1.979641 78.460718 21.274175 153.352504 49.435271 225.846415 11.766319 30.335914 37.167071 44.416462 69.510508 43.858816 38.059303-0.641292 76.118607-1.84023 114.094263-4.042929a316.77051 316.77051 0 0 0 47.985393-7.751272c22.473112-4.851516 38.338126-17.28701 44.611637-40.680237 3.262226-12.045142 8.894445-23.448992 12.351847-35.466252 2.509405-8.727152 7.556096-12.073024 16.06019-14.582429 15.363133-4.489046 32.901083-7.779154 44.611638-17.565833 19.517591-16.56207 35.549899-37.585305 52.61385-57.102896 5.576455-6.329276 5.046692-13.299844-3.206462-17.203363-19.517591-9.312679-39.035183-18.681123-59.249831-26.7391-7.10998-2.788227-8.978092-5.297632-7.946448-12.853728 1.868112-13.941137 2.119053-27.882274 2.955521-40.457179-129.26222 29.220623-255.708331 26.432395-382.851498-1.087409zM292.093467 789.514457l-12.547023-10.818322c-1.115291-6.580217-1.951759-11.571144-3.011285-17.872537l6.329276-4.098695-0.97588-3.178579-20.019472 2.788228-12.714317-7.583979c-0.278823-4.712104-0.61341-10.037618-0.752821-12.602787l11.431732-11.626908L240.790084 716.602312l-14.610311-14.693958c0-0.808586 0.306705-4.015047 0.724939-9.675149a42.631996 42.631996 0 0 0-8.141624 5.827395c-0.947997 1.198938-0.557645 3.596813-0.473999 5.409161 2.788227 56.65678 31.925203 108.936043 99.0936 117.105549 18.402301 2.258464 36.91613 3.708342 55.402078 5.018809 8.978092 0.641292 18.011949 0 26.069926 0-10.734675-58.190305-21.21841-114.930731-31.674263-171.69904l-3.513167-0.641293c-1.449878 13.745961-2.788227 27.491922-4.461163 42.18588-10.734675-2.788227-9.284797 4.572693-10.121266 9.619385l-11.152909 8.950209 1.254702 1.366232-28.161096 7.918566 22.640406 13.271962c2.788227 4.265988 5.409161 8.615623 7.695508 12.2682 0.473999 5.102456 0.97588 10.232794 1.254702 13.076786l-3.345873 16.366895-7.918566 11.152909-13.941136 7.807037-12.770082-1.115291z m64.686875-169.050224c0 5.409161-0.278823 8.894445 0 12.296082a23.42111 23.42111 0 0 0 2.230582 8.364682 74.752375 74.752375 0 0 0 7.890683 10.009737c0-13.718079-0.557645-22.947111 0.223058-32.064615 0.36247-4.154459 2.314229-10.121265 5.381279-11.766319 20.381942-10.901969 41.82341-18.123478 65.467578-12.574906 8.58774 2.007524 17.28701 3.485284 25.87475 5.576455 11.905731 2.788227 17.314892-2.565169 15.391015-13.941137-4.600575-27.408275-9.368444-54.844432-15.418897-81.946002-2.788227-12.714317-8.727152-24.759459-13.24408-37.083423a15.44678 15.44678 0 0 0-5.576455 10.651028 62.930291 62.930291 0 0 1-22.919229 44.611638 327.477303 327.477303 0 0 1-33.458728 25.094046C370.163833 559.374171 350.646242 570.248258 329.399949 582.767399l22.919229 27.882273c-5.687984 5.353397-3.903518 9.312679 4.461164 9.814561z m-122.096476 75.588843c18.653241 21.302057 58.273952 29.443681 81.527768 17.426421 17.203363-8.894445 31.03297-21.21841 34.183667-41.321529 3.373755-21.58088 0.697057-42.520467-10.706793-61.870765-13.718079-23.337463-18.346536-24.620048-40.680237-10.149148-3.513166 2.258464-7.193627 4.321752-10.539499 6.803275-9.173268 6.775392-6.886922 19.768532 2.509404 25.595927 18.207125 11.152909 31.311793 1.505643 44.834696-8.615622 0.947997-0.724939 1.979641-1.310467 4.210223-2.788228l2.983404 10.901969c-14.917016 9.870325-33.793316 7.72339-42.631997 27.631333-9.479973 21.329939 4.739986 32.454966 14.526665 47.818099l-23.198052 7.305156c0.947997-8.699269 3.011286-15.614073 2.035406-22.082761s-3.06705-16.31113-7.862801-19.043592c-19.517591-11.152909-23.67205-9.535738-39.258241 8.002212-3.987165 4.516928-7.667625 9.256915-11.933613 14.387253zM475.168475 632.955491c60.058417 10.957733 120.116834 10.678911 180.175252 4.516929V632.955491z m-188.874521 37.250718c4.377517-7.807037 8.197388-12.240318 9.061739-17.175481 0.390352-2.258464-6.886922-8.364682-7.583978-7.890683-4.516928 2.788227-9.507855 6.608099-11.543261 11.152909-0.86435 2.119053 4.851516 7.054215 10.0655 13.913255z m87.633986-543.704334l-3.317991-4.238106L353.434469 133.360914l16.394777 11.375968c1.868112-8.448329 3.122815-13.271962 4.098694-18.123478z m91.73268 5.938924l-0.697057 5.548573 19.266651 8.113741v-17.593714z m-81.806591-9.396326c-2.063288 9.730913-3.06705 14.331489-5.046691 23.67205l18.848417-9.926089z m242.018135 471.963244l-2.927639 5.26975c2.230582 9.870325 8.364682 11.320203 16.868775 8.030095 0.808586-1.505643 1.58929-3.011286 2.369994-4.516929z m-38.756361 20.911705l-16.199601-17.78889-3.541048 3.429519c1.031644 9.089621 3.819871 16.450541 19.740649 14.4709z" p-id="6749"></path><path d="M616.50372 702.019883a30.670501 30.670501 0 0 1-1.868113 6.078335c-6.078336 10.762558-11.375968 20.493471 8.364682 22.305819 3.457402 0.306705 8.58774 7.611861 8.978093 12.045142 1.923877 21.246292 2.788227 42.604114 3.290108 63.934054 0.223058 10.79044-5.576455 17.203363-17.203363 17.426421q-54.258904 1.087409-108.517809 2.425757c-8.699269 0.195176-13.021022-4.377517-13.216197-12.63067-0.557645-22.724053-0.836468-45.448106-1.143173-68.172158 0-9.312679 3.736225-14.136313 13.941136-15.195839 20.632882-2.146935 20.577118-2.620934 13.271963-21.803938a63.209114 63.209114 0 0 1-2.258465-6.580217 27.073688 27.073688 0 0 1 1.22682-6.078335c10.372206 20.158884 20.326177 34.044256 45.754811 32.62226 22.668288-1.282585 38.310244-6.608099 46.423986-30.670501z m-51.665853 114.651909c16.227483 0 32.454966-0.306705 48.654567 0 10.567382 0.278823 15.195839-3.652578 14.861252-14.638194q-0.752821-25.735338 0.25094-51.470677c0.418234-10.093383-4.265988-13.160433-13.299844-12.965257-33.319317 0.669175-66.638634 1.338349-99.957951 1.756583-8.615623 0-12.853728 3.568931-12.714316 12.463376q0.36247 25.735338 0.25094 51.442795c0 10.037618 4.65634 13.941137 14.666076 13.522903 15.753485-0.501881 31.534851-0.111529 47.288336-0.111529zM725.049411 780.731541c7.751272-28.216861 15.44678-56.154899 22.724052-82.53153 8.95021 3.541049 18.179242 7.221509 27.436158 10.846205 29.276387 11.487497 29.973444 14.219959 10.260676 39.230359-18.876299 24.090284-36.330602 33.59814-60.420886 32.454966z" p-id="6750"></path></svg>